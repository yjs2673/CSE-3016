`timescale 1ns / 1ps

module convert_tb;
reg a, b, c, d;
wire e, f, g, h;

convert u_convert (
   .a(a ),
   .b(b ),
   .c(c ),
   .d(d ),
   .e(e ),
   .f(f ),
   .g(g ),
   .h(h )
);

initial begin
   a = 1'b0;
   b = 1'b0;
   c = 1'b0;
   d = 1'b0;
end

always@(a or b or c or d) begin
   a <= #50 ~a;
   b <= #100 ~b;
   c <= #150 ~c;
   d <= #200 ~d;
end

initial begin
   #1000
   $finish;
end

endmodule
